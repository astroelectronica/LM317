.title KiCad schematic
.include "C:/AE/LM317/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/LM317/_models/C3216X7R2A105M160AA_p.mod"
.include "C:/AE/LM317/_models/LM317.lib"
R1 /ADJ /VOUT {RADJ}
XU3 /VOUT 0 C3216X7R2A105M160AA_p
XU2 /VIN 0 C2012X7R2A104K125AA_p
XU1 /VIN /ADJ /VOUT LM317
R2 /ADJ 0 {RREF}
V1 /VIN 0 {VSOURCE}
I1 /VOUT 0 {ILOAD}
.end
